-- megafunction wizard: %Flash Memory%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altufm_parallel 

-- ============================================================
-- File Name: flash.vhd
-- Megafunction Name(s):
-- 			altufm_parallel
--
-- Simulation Library Files(s):
-- 			lpm;maxii
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.1 Build 304 01/25/2010 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2010 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altufm_parallel ACCESS_MODE="READ_WRITE" CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="MAX II" ERASE_TIME=500000000 LPM_FILE="tstdata.mif" OSC_FREQUENCY=180000 PROGRAM_TIME=1600000 WIDTH_ADDRESS=9 WIDTH_DATA=8 WIDTH_UFM_ADDRESS=9 addr data_valid datain dataout nbusy nerase nread nwrite
--VERSION_BEGIN 9.1SP1 cbx_a_gray2bin 2010:01:25:21:24:34:SJ cbx_a_graycounter 2010:01:25:21:24:34:SJ cbx_altufm_parallel 2010:01:25:21:24:34:SJ cbx_cycloneii 2010:01:25:21:24:34:SJ cbx_lpm_add_sub 2010:01:25:21:24:34:SJ cbx_lpm_compare 2010:01:25:21:24:34:SJ cbx_lpm_counter 2010:01:25:21:24:34:SJ cbx_lpm_decode 2010:01:25:21:24:34:SJ cbx_lpm_mux 2010:01:25:21:24:34:SJ cbx_maxii 2010:01:25:21:24:34:SJ cbx_mgl 2010:01:25:21:38:39:SJ cbx_stratix 2010:01:25:21:24:34:SJ cbx_stratixii 2010:01:25:21:24:34:SJ cbx_util_mgl 2010:01:25:21:24:34:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

 LIBRARY maxii;
 USE maxii.all;

--synthesis_resources = lpm_counter 1 lut 71 maxii_ufm 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  flash_altufm_parallel_22p IS 
	 PORT 
	 ( 
		 addr	:	IN  STD_LOGIC_VECTOR (8 DOWNTO 0);
		 data_valid	:	OUT  STD_LOGIC;
		 datain	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 dataout	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 nbusy	:	OUT  STD_LOGIC;
		 nerase	:	IN  STD_LOGIC := '1';
		 nread	:	IN  STD_LOGIC;
		 nwrite	:	IN  STD_LOGIC := '1'
	 ); 
 END flash_altufm_parallel_22p;

 ARCHITECTURE RTL OF flash_altufm_parallel_22p IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "suppress_da_rule_internal=c101;suppress_da_rule_internal=c103;suppress_da_rule_internal=c104;suppress_da_rule_internal=r101;suppress_da_rule_internal=s104;suppress_da_rule_internal=s102";

	 SIGNAL	 A	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 data_valid_out_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 data_valid_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_data_valid_reg_w_lg_q100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 deco1_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 deco2_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 deco3_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 decode_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 gated_clk1_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 gated_clk2_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 piso_sipo_dffe	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 program_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_program_dffe_clrn	:	STD_LOGIC;
	 SIGNAL	 real_decode2_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_real_decode2_dffe_w_lg_q27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 real_decode_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_tmp_do_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 tmp_do	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_tmp_do_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL  wire_cntr2_cnt_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_ufm_program45w46w47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cntr2_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_maxii_ufm_block1_bgpbusy	:	STD_LOGIC;
	 SIGNAL  wire_maxii_ufm_block1_busy	:	STD_LOGIC;
	 SIGNAL  wire_maxii_ufm_block1_drdout	:	STD_LOGIC;
	 SIGNAL  wire_maxii_ufm_block1_osc	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_q363w72w73w74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_mux_nread20w21w22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_q363w72w73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_tmp_read36w37w38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_mux_nread18w19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_tmp_read34w35w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_control_mux7w12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_control_mux7w8w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_control_mux7w10w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_mux_nread20w21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_q253w62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_q363w72w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_q363w127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_q363w126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_q363w128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_q43w54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_op110w114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_op110w117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_op110w111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_tmp_read36w37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_addr144w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_mux_nread18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_q160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_q3124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_q475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_q481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_q466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shiftin143w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_tmp_read34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_ufm_drdout160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_piso_sipo_q_range166w171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_piso_sipo_q_range266w271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_piso_sipo_q_range276w281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_piso_sipo_q_range286w291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_piso_sipo_q_range296w301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_piso_sipo_q_range306w311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_piso_sipo_q_range176w181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_piso_sipo_q_range186w191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_piso_sipo_q_range196w201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_piso_sipo_q_range206w211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_piso_sipo_q_range216w221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_piso_sipo_q_range226w231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_piso_sipo_q_range236w241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_piso_sipo_q_range246w251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_piso_sipo_q_range256w261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tmp_di_range156w158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tmp_di_range258w260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tmp_di_range268w270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tmp_di_range278w280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tmp_di_range288w290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tmp_di_range298w300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tmp_di_range308w310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tmp_di_range168w170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tmp_di_range178w180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tmp_di_range188w190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tmp_di_range198w200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tmp_di_range208w210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tmp_di_range218w220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tmp_di_range228w230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tmp_di_range238w240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tmp_di_range248w250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_add_load142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_control_mux7w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_data_load159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dly_tmp_decode41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_mux_nerase14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_mux_nread20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_mux_nwrite17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_q059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_q161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_q253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_q363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_q43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_op110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_tmp_decode99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_tmp_erase30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_tmp_read36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_tmp_write33w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_ufm_bgpbusy25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_ufm_osc321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_ufm_drdout160w161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_piso_sipo_q_range166w171w172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_piso_sipo_q_range266w271w272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_piso_sipo_q_range276w281w282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_piso_sipo_q_range286w291w292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_piso_sipo_q_range296w301w302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_piso_sipo_q_range306w311w312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_piso_sipo_q_range176w181w182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_piso_sipo_q_range186w191w192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_piso_sipo_q_range196w201w202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_piso_sipo_q_range206w211w212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_piso_sipo_q_range216w221w222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_piso_sipo_q_range226w231w232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_piso_sipo_q_range236w241w242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_piso_sipo_q_range246w251w252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_piso_sipo_q_range256w261w262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_q363w64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_q363w64w65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_q31w2w76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_q31w2w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_q31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  add_en :	STD_LOGIC;
	 SIGNAL  add_load :	STD_LOGIC;
	 SIGNAL  arclk :	STD_LOGIC;
	 SIGNAL  busy_arclk :	STD_LOGIC;
	 SIGNAL  busy_drclk :	STD_LOGIC;
	 SIGNAL  control_mux :	STD_LOGIC;
	 SIGNAL  copy_tmp_decode :	STD_LOGIC;
	 SIGNAL  data_en :	STD_LOGIC;
	 SIGNAL  data_load :	STD_LOGIC;
	 SIGNAL  data_valid_en :	STD_LOGIC;
	 SIGNAL  dly_tmp_decode :	STD_LOGIC;
	 SIGNAL  drclk :	STD_LOGIC;
	 SIGNAL  drshft :	STD_LOGIC;
	 SIGNAL  erase :	STD_LOGIC;
	 SIGNAL  erase_op :	STD_LOGIC;
	 SIGNAL  gated1 :	STD_LOGIC;
	 SIGNAL  gated2 :	STD_LOGIC;
	 SIGNAL  hold_decode :	STD_LOGIC;
	 SIGNAL  in_erase :	STD_LOGIC;
	 SIGNAL  in_program :	STD_LOGIC;
	 SIGNAL  in_read_data_en :	STD_LOGIC;
	 SIGNAL  in_read_drclk :	STD_LOGIC;
	 SIGNAL  in_read_drshft :	STD_LOGIC;
	 SIGNAL  in_write_data_en :	STD_LOGIC;
	 SIGNAL  in_write_data_load :	STD_LOGIC;
	 SIGNAL  in_write_drclk :	STD_LOGIC;
	 SIGNAL  in_write_drshft :	STD_LOGIC;
	 SIGNAL  mux_nerase :	STD_LOGIC;
	 SIGNAL  mux_nread :	STD_LOGIC;
	 SIGNAL  mux_nwrite :	STD_LOGIC;
	 SIGNAL  oscena	:	STD_LOGIC;
	 SIGNAL  piso_sipo_d :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  piso_sipo_q :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  program1 :	STD_LOGIC;
	 SIGNAL  q0 :	STD_LOGIC;
	 SIGNAL  q1 :	STD_LOGIC;
	 SIGNAL  q2 :	STD_LOGIC;
	 SIGNAL  q3 :	STD_LOGIC;
	 SIGNAL  q4 :	STD_LOGIC;
	 SIGNAL  read_data_en :	STD_LOGIC;
	 SIGNAL  read_drclk :	STD_LOGIC;
	 SIGNAL  read_drshft :	STD_LOGIC;
	 SIGNAL  read_op :	STD_LOGIC;
	 SIGNAL  real_decode :	STD_LOGIC;
	 SIGNAL  shiftin :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  start_decode :	STD_LOGIC;
	 SIGNAL  start_op :	STD_LOGIC;
	 SIGNAL  stop_op :	STD_LOGIC;
	 SIGNAL  tmp_add_en :	STD_LOGIC;
	 SIGNAL  tmp_add_load :	STD_LOGIC;
	 SIGNAL  tmp_arclk :	STD_LOGIC;
	 SIGNAL  tmp_arclk0 :	STD_LOGIC;
	 SIGNAL  tmp_ardin :	STD_LOGIC;
	 SIGNAL  tmp_arshft :	STD_LOGIC;
	 SIGNAL  tmp_data_valid2 :	STD_LOGIC;
	 SIGNAL  tmp_decode :	STD_LOGIC;
	 SIGNAL  tmp_di :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  tmp_drclk :	STD_LOGIC;
	 SIGNAL  tmp_drdin :	STD_LOGIC;
	 SIGNAL  tmp_erase :	STD_LOGIC;
	 SIGNAL  tmp_read :	STD_LOGIC;
	 SIGNAL  tmp_write :	STD_LOGIC;
	 SIGNAL  ufm_arclk :	STD_LOGIC;
	 SIGNAL  ufm_ardin :	STD_LOGIC;
	 SIGNAL  ufm_arshft :	STD_LOGIC;
	 SIGNAL  ufm_bgpbusy :	STD_LOGIC;
	 SIGNAL  ufm_busy :	STD_LOGIC;
	 SIGNAL  ufm_drclk :	STD_LOGIC;
	 SIGNAL  ufm_drdin :	STD_LOGIC;
	 SIGNAL  ufm_drdout :	STD_LOGIC;
	 SIGNAL  ufm_drshft :	STD_LOGIC;
	 SIGNAL  ufm_erase :	STD_LOGIC;
	 SIGNAL  ufm_osc :	STD_LOGIC;
	 SIGNAL  ufm_oscena :	STD_LOGIC;
	 SIGNAL  ufm_program :	STD_LOGIC;
	 SIGNAL  write_data_en :	STD_LOGIC;
	 SIGNAL  write_data_load :	STD_LOGIC;
	 SIGNAL  write_drclk :	STD_LOGIC;
	 SIGNAL  write_drshft :	STD_LOGIC;
	 SIGNAL  write_op :	STD_LOGIC;
	 SIGNAL  X_var :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  Y_var :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  Z_var :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_piso_sipo_q_range166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_piso_sipo_q_range266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_piso_sipo_q_range276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_piso_sipo_q_range286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_piso_sipo_q_range296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_piso_sipo_q_range306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_piso_sipo_q_range176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_piso_sipo_q_range186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_piso_sipo_q_range196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_piso_sipo_q_range206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_piso_sipo_q_range216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_piso_sipo_q_range226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_piso_sipo_q_range236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_piso_sipo_q_range246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_piso_sipo_q_range256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tmp_di_range156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tmp_di_range258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tmp_di_range268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tmp_di_range278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tmp_di_range288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tmp_di_range298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tmp_di_range308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tmp_di_range168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tmp_di_range178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tmp_di_range188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tmp_di_range198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tmp_di_range208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tmp_di_range218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tmp_di_range228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tmp_di_range238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tmp_di_range248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  maxii_ufm
	 GENERIC 
	 (
		ADDRESS_WIDTH	:	NATURAL := 9;
		ERASE_TIME	:	NATURAL := 500000000;
		INIT_FILE	:	STRING := "UNUSED";
		mem1	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem10	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem11	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem12	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem13	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem14	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem15	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem16	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem2	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem3	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem4	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem5	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem6	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem7	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem8	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem9	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		OSC_SIM_SETTING	:	NATURAL := 180000;
		PROGRAM_TIME	:	NATURAL := 1600000;
		lpm_type	:	STRING := "maxii_ufm"
	 );
	 PORT
	 ( 
		arclk	:	IN STD_LOGIC := '0';
		ardin	:	IN STD_LOGIC := '0';
		arshft	:	IN STD_LOGIC := '1';
		bgpbusy	:	OUT STD_LOGIC;
		busy	:	OUT STD_LOGIC;
		drclk	:	IN STD_LOGIC := '0';
		drdin	:	IN STD_LOGIC := '0';
		drdout	:	OUT STD_LOGIC;
		drshft	:	IN STD_LOGIC := '1';
		erase	:	IN STD_LOGIC := '0';
		osc	:	OUT STD_LOGIC;
		oscena	:	IN STD_LOGIC := '0';
		program	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w_lg_w_lg_w_lg_q363w72w73w74w(0) <= wire_w_lg_w_lg_w_lg_q363w72w73w(0) AND wire_w_lg_q059w(0);
	wire_w_lg_w_lg_w_lg_mux_nread20w21w22w(0) <= wire_w_lg_w_lg_mux_nread20w21w(0) AND mux_nerase;
	wire_w_lg_w_lg_w_lg_q363w72w73w(0) <= wire_w_lg_w_lg_q363w72w(0) AND wire_w_lg_q161w(0);
	wire_w_lg_w_lg_w_lg_tmp_read36w37w38w(0) <= wire_w_lg_w_lg_tmp_read36w37w(0) AND tmp_erase;
	wire_w_lg_w_lg_mux_nread18w19w(0) <= wire_w_lg_mux_nread18w(0) AND mux_nerase;
	wire_w_lg_w_lg_tmp_read34w35w(0) <= wire_w_lg_tmp_read34w(0) AND tmp_erase;
	wire_w_lg_w_lg_control_mux7w12w(0) <= wire_w_lg_control_mux7w(0) AND nerase;
	wire_w_lg_w_lg_control_mux7w8w(0) <= wire_w_lg_control_mux7w(0) AND nread;
	wire_w_lg_w_lg_control_mux7w10w(0) <= wire_w_lg_control_mux7w(0) AND nwrite;
	wire_w_lg_w_lg_mux_nread20w21w(0) <= wire_w_lg_mux_nread20w(0) AND mux_nwrite;
	wire_w_lg_w_lg_q253w62w(0) <= wire_w_lg_q253w(0) AND wire_w_lg_q161w(0);
	wire_w_lg_w_lg_q363w72w(0) <= wire_w_lg_q363w(0) AND wire_w_lg_q253w(0);
	wire_w_lg_w_lg_q363w127w(0) <= wire_w_lg_q363w(0) AND q0;
	wire_w_lg_w_lg_q363w126w(0) <= wire_w_lg_q363w(0) AND q1;
	wire_w_lg_w_lg_q363w128w(0) <= wire_w_lg_q363w(0) AND q2;
	wire_w_lg_w_lg_q43w54w(0) <= wire_w_lg_q43w(0) AND q3;
	wire_w_lg_w_lg_read_op110w114w(0) <= wire_w_lg_read_op110w(0) AND write_data_en;
	wire_w_lg_w_lg_read_op110w117w(0) <= wire_w_lg_read_op110w(0) AND write_drclk;
	wire_w_lg_w_lg_read_op110w111w(0) <= wire_w_lg_read_op110w(0) AND write_drshft;
	wire_w_lg_w_lg_tmp_read36w37w(0) <= wire_w_lg_tmp_read36w(0) AND tmp_write;
	loop0 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_addr144w(i) <= addr(i) AND add_load;
	END GENERATE loop0;
	wire_w_lg_mux_nread18w(0) <= mux_nread AND wire_w_lg_mux_nwrite17w(0);
	wire_w_lg_q160w(0) <= q1 AND wire_w_lg_q059w(0);
	wire_w_lg_q3124w(0) <= q3 AND wire_w_lg_q253w(0);
	wire_w_lg_q475w(0) <= q4 AND wire_w_lg_w_lg_w_lg_w_lg_q363w72w73w74w(0);
	wire_w_lg_q481w(0) <= q4 AND wire_w_lg_q363w(0);
	wire_w_lg_q466w(0) <= q4 AND wire_w_lg_w_lg_w_lg_q363w64w65w(0);
	loop1 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_shiftin143w(i) <= shiftin(i) AND wire_w_lg_add_load142w(0);
	END GENERATE loop1;
	wire_w_lg_tmp_read34w(0) <= tmp_read AND wire_w_lg_tmp_write33w(0);
	wire_w_lg_ufm_drdout160w(0) <= ufm_drdout AND wire_w_lg_data_load159w(0);
	wire_w_lg_w_piso_sipo_q_range166w171w(0) <= wire_w_piso_sipo_q_range166w(0) AND wire_w_lg_data_load159w(0);
	wire_w_lg_w_piso_sipo_q_range266w271w(0) <= wire_w_piso_sipo_q_range266w(0) AND wire_w_lg_data_load159w(0);
	wire_w_lg_w_piso_sipo_q_range276w281w(0) <= wire_w_piso_sipo_q_range276w(0) AND wire_w_lg_data_load159w(0);
	wire_w_lg_w_piso_sipo_q_range286w291w(0) <= wire_w_piso_sipo_q_range286w(0) AND wire_w_lg_data_load159w(0);
	wire_w_lg_w_piso_sipo_q_range296w301w(0) <= wire_w_piso_sipo_q_range296w(0) AND wire_w_lg_data_load159w(0);
	wire_w_lg_w_piso_sipo_q_range306w311w(0) <= wire_w_piso_sipo_q_range306w(0) AND wire_w_lg_data_load159w(0);
	wire_w_lg_w_piso_sipo_q_range176w181w(0) <= wire_w_piso_sipo_q_range176w(0) AND wire_w_lg_data_load159w(0);
	wire_w_lg_w_piso_sipo_q_range186w191w(0) <= wire_w_piso_sipo_q_range186w(0) AND wire_w_lg_data_load159w(0);
	wire_w_lg_w_piso_sipo_q_range196w201w(0) <= wire_w_piso_sipo_q_range196w(0) AND wire_w_lg_data_load159w(0);
	wire_w_lg_w_piso_sipo_q_range206w211w(0) <= wire_w_piso_sipo_q_range206w(0) AND wire_w_lg_data_load159w(0);
	wire_w_lg_w_piso_sipo_q_range216w221w(0) <= wire_w_piso_sipo_q_range216w(0) AND wire_w_lg_data_load159w(0);
	wire_w_lg_w_piso_sipo_q_range226w231w(0) <= wire_w_piso_sipo_q_range226w(0) AND wire_w_lg_data_load159w(0);
	wire_w_lg_w_piso_sipo_q_range236w241w(0) <= wire_w_piso_sipo_q_range236w(0) AND wire_w_lg_data_load159w(0);
	wire_w_lg_w_piso_sipo_q_range246w251w(0) <= wire_w_piso_sipo_q_range246w(0) AND wire_w_lg_data_load159w(0);
	wire_w_lg_w_piso_sipo_q_range256w261w(0) <= wire_w_piso_sipo_q_range256w(0) AND wire_w_lg_data_load159w(0);
	wire_w_lg_w_tmp_di_range156w158w(0) <= wire_w_tmp_di_range156w(0) AND data_load;
	wire_w_lg_w_tmp_di_range258w260w(0) <= wire_w_tmp_di_range258w(0) AND data_load;
	wire_w_lg_w_tmp_di_range268w270w(0) <= wire_w_tmp_di_range268w(0) AND data_load;
	wire_w_lg_w_tmp_di_range278w280w(0) <= wire_w_tmp_di_range278w(0) AND data_load;
	wire_w_lg_w_tmp_di_range288w290w(0) <= wire_w_tmp_di_range288w(0) AND data_load;
	wire_w_lg_w_tmp_di_range298w300w(0) <= wire_w_tmp_di_range298w(0) AND data_load;
	wire_w_lg_w_tmp_di_range308w310w(0) <= wire_w_tmp_di_range308w(0) AND data_load;
	wire_w_lg_w_tmp_di_range168w170w(0) <= wire_w_tmp_di_range168w(0) AND data_load;
	wire_w_lg_w_tmp_di_range178w180w(0) <= wire_w_tmp_di_range178w(0) AND data_load;
	wire_w_lg_w_tmp_di_range188w190w(0) <= wire_w_tmp_di_range188w(0) AND data_load;
	wire_w_lg_w_tmp_di_range198w200w(0) <= wire_w_tmp_di_range198w(0) AND data_load;
	wire_w_lg_w_tmp_di_range208w210w(0) <= wire_w_tmp_di_range208w(0) AND data_load;
	wire_w_lg_w_tmp_di_range218w220w(0) <= wire_w_tmp_di_range218w(0) AND data_load;
	wire_w_lg_w_tmp_di_range228w230w(0) <= wire_w_tmp_di_range228w(0) AND data_load;
	wire_w_lg_w_tmp_di_range238w240w(0) <= wire_w_tmp_di_range238w(0) AND data_load;
	wire_w_lg_w_tmp_di_range248w250w(0) <= wire_w_tmp_di_range248w(0) AND data_load;
	wire_w_lg_add_load142w(0) <= NOT add_load;
	wire_w_lg_control_mux7w(0) <= NOT control_mux;
	wire_w_lg_data_load159w(0) <= NOT data_load;
	wire_w_lg_dly_tmp_decode41w(0) <= NOT dly_tmp_decode;
	wire_w_lg_mux_nerase14w(0) <= NOT mux_nerase;
	wire_w_lg_mux_nread20w(0) <= NOT mux_nread;
	wire_w_lg_mux_nwrite17w(0) <= NOT mux_nwrite;
	wire_w_lg_q059w(0) <= NOT q0;
	wire_w_lg_q161w(0) <= NOT q1;
	wire_w_lg_q253w(0) <= NOT q2;
	wire_w_lg_q363w(0) <= NOT q3;
	wire_w_lg_q43w(0) <= NOT q4;
	wire_w_lg_read_op110w(0) <= NOT read_op;
	wire_w_lg_tmp_decode99w(0) <= NOT tmp_decode;
	wire_w_lg_tmp_erase30w(0) <= NOT tmp_erase;
	wire_w_lg_tmp_read36w(0) <= NOT tmp_read;
	wire_w_lg_tmp_write33w(0) <= NOT tmp_write;
	wire_w_lg_ufm_bgpbusy25w(0) <= NOT ufm_bgpbusy;
	wire_w_lg_ufm_osc321w(0) <= NOT ufm_osc;
	wire_w_lg_w_lg_ufm_drdout160w161w(0) <= wire_w_lg_ufm_drdout160w(0) OR wire_w_lg_w_tmp_di_range156w158w(0);
	wire_w_lg_w_lg_w_piso_sipo_q_range166w171w172w(0) <= wire_w_lg_w_piso_sipo_q_range166w171w(0) OR wire_w_lg_w_tmp_di_range168w170w(0);
	wire_w_lg_w_lg_w_piso_sipo_q_range266w271w272w(0) <= wire_w_lg_w_piso_sipo_q_range266w271w(0) OR wire_w_lg_w_tmp_di_range268w270w(0);
	wire_w_lg_w_lg_w_piso_sipo_q_range276w281w282w(0) <= wire_w_lg_w_piso_sipo_q_range276w281w(0) OR wire_w_lg_w_tmp_di_range278w280w(0);
	wire_w_lg_w_lg_w_piso_sipo_q_range286w291w292w(0) <= wire_w_lg_w_piso_sipo_q_range286w291w(0) OR wire_w_lg_w_tmp_di_range288w290w(0);
	wire_w_lg_w_lg_w_piso_sipo_q_range296w301w302w(0) <= wire_w_lg_w_piso_sipo_q_range296w301w(0) OR wire_w_lg_w_tmp_di_range298w300w(0);
	wire_w_lg_w_lg_w_piso_sipo_q_range306w311w312w(0) <= wire_w_lg_w_piso_sipo_q_range306w311w(0) OR wire_w_lg_w_tmp_di_range308w310w(0);
	wire_w_lg_w_lg_w_piso_sipo_q_range176w181w182w(0) <= wire_w_lg_w_piso_sipo_q_range176w181w(0) OR wire_w_lg_w_tmp_di_range178w180w(0);
	wire_w_lg_w_lg_w_piso_sipo_q_range186w191w192w(0) <= wire_w_lg_w_piso_sipo_q_range186w191w(0) OR wire_w_lg_w_tmp_di_range188w190w(0);
	wire_w_lg_w_lg_w_piso_sipo_q_range196w201w202w(0) <= wire_w_lg_w_piso_sipo_q_range196w201w(0) OR wire_w_lg_w_tmp_di_range198w200w(0);
	wire_w_lg_w_lg_w_piso_sipo_q_range206w211w212w(0) <= wire_w_lg_w_piso_sipo_q_range206w211w(0) OR wire_w_lg_w_tmp_di_range208w210w(0);
	wire_w_lg_w_lg_w_piso_sipo_q_range216w221w222w(0) <= wire_w_lg_w_piso_sipo_q_range216w221w(0) OR wire_w_lg_w_tmp_di_range218w220w(0);
	wire_w_lg_w_lg_w_piso_sipo_q_range226w231w232w(0) <= wire_w_lg_w_piso_sipo_q_range226w231w(0) OR wire_w_lg_w_tmp_di_range228w230w(0);
	wire_w_lg_w_lg_w_piso_sipo_q_range236w241w242w(0) <= wire_w_lg_w_piso_sipo_q_range236w241w(0) OR wire_w_lg_w_tmp_di_range238w240w(0);
	wire_w_lg_w_lg_w_piso_sipo_q_range246w251w252w(0) <= wire_w_lg_w_piso_sipo_q_range246w251w(0) OR wire_w_lg_w_tmp_di_range248w250w(0);
	wire_w_lg_w_lg_w_piso_sipo_q_range256w261w262w(0) <= wire_w_lg_w_piso_sipo_q_range256w261w(0) OR wire_w_lg_w_tmp_di_range258w260w(0);
	wire_w_lg_w_lg_q363w64w(0) <= wire_w_lg_q363w(0) OR wire_w_lg_w_lg_q253w62w(0);
	wire_w_lg_w_lg_w_lg_q363w64w65w(0) <= wire_w_lg_w_lg_q363w64w(0) OR wire_w_lg_q160w(0);
	wire_w_lg_w_lg_w_lg_q31w2w76w(0) <= wire_w_lg_w_lg_q31w2w(0) OR q0;
	wire_w_lg_w_lg_q31w2w(0) <= wire_w_lg_q31w(0) OR q1;
	wire_w_lg_q31w(0) <= q3 OR q2;
	add_en <= (tmp_add_en AND ((read_op OR write_op) OR erase_op));
	add_load <= (tmp_add_load AND ((read_op OR write_op) OR erase_op));
	arclk <= (tmp_arclk0 AND ((read_op OR write_op) OR erase_op));
	busy_arclk <= arclk;
	busy_drclk <= drclk;
	control_mux <= ((wire_w_lg_q43w(0) AND wire_w_lg_w_lg_q31w2w(0)) OR q4);
	copy_tmp_decode <= tmp_decode;
	data_en <= (wire_w_lg_w_lg_read_op110w114w(0) OR (read_op AND read_data_en));
	data_load <= (write_data_load AND write_op);
	data_valid <= data_valid_out_reg;
	data_valid_en <= ((q4 AND q3) AND q1);
	dataout <= tmp_do;
	dly_tmp_decode <= decode_dffe;
	drclk <= (wire_w_lg_w_lg_read_op110w117w(0) OR (read_op AND read_drclk));
	drshft <= (wire_w_lg_w_lg_read_op110w111w(0) OR (read_op AND read_drshft));
	erase <= (in_erase AND erase_op);
	erase_op <= ((tmp_read AND tmp_write) AND wire_w_lg_tmp_erase30w(0));
	gated1 <= gated_clk1_dffe;
	gated2 <= gated_clk2_dffe;
	hold_decode <= (wire_real_decode2_dffe_w_lg_q27w(0) AND real_decode);
	in_erase <= (((wire_w_lg_w_lg_q43w54w(0) AND wire_w_lg_q253w(0)) AND q1) AND q0);
	in_program <= (((wire_w_lg_q481w(0) AND wire_w_lg_q253w(0)) AND wire_w_lg_q161w(0)) AND q0);
	in_read_data_en <= ((wire_w_lg_q43w(0) AND ((q3 AND q2) OR (q3 AND q1))) OR wire_w_lg_q466w(0));
	in_read_drclk <= ((wire_w_lg_q43w(0) AND ((q3 AND q2) OR (q3 AND q1))) OR wire_w_lg_q466w(0));
	in_read_drshft <= (NOT (((wire_w_lg_w_lg_q43w54w(0) AND wire_w_lg_q253w(0)) AND q1) AND q0));
	in_write_data_en <= (wire_w_lg_q43w(0) OR wire_w_lg_w_lg_w_lg_w_lg_q363w72w73w74w(0));
	in_write_data_load <= (NOT ((wire_w_lg_q43w(0) AND wire_w_lg_w_lg_w_lg_q31w2w76w(0)) OR wire_w_lg_q475w(0)));
	in_write_drclk <= wire_w_lg_q43w(0);
	in_write_drshft <= in_write_data_en;
	mux_nerase <= (wire_w_lg_w_lg_control_mux7w12w(0) OR (control_mux AND data_valid_en));
	mux_nread <= (wire_w_lg_w_lg_control_mux7w8w(0) OR (control_mux AND data_valid_en));
	mux_nwrite <= (wire_w_lg_w_lg_control_mux7w10w(0) OR (control_mux AND data_valid_en));
	nbusy <= (wire_w_lg_dly_tmp_decode41w(0) AND wire_w_lg_ufm_bgpbusy25w(0));
	oscena <= '1';
	piso_sipo_d <= ( wire_w_lg_w_lg_w_piso_sipo_q_range306w311w312w & wire_w_lg_w_lg_w_piso_sipo_q_range296w301w302w & wire_w_lg_w_lg_w_piso_sipo_q_range286w291w292w & wire_w_lg_w_lg_w_piso_sipo_q_range276w281w282w & wire_w_lg_w_lg_w_piso_sipo_q_range266w271w272w & wire_w_lg_w_lg_w_piso_sipo_q_range256w261w262w & wire_w_lg_w_lg_w_piso_sipo_q_range246w251w252w & wire_w_lg_w_lg_w_piso_sipo_q_range236w241w242w & wire_w_lg_w_lg_w_piso_sipo_q_range226w231w232w & wire_w_lg_w_lg_w_piso_sipo_q_range216w221w222w & wire_w_lg_w_lg_w_piso_sipo_q_range206w211w212w & wire_w_lg_w_lg_w_piso_sipo_q_range196w201w202w & wire_w_lg_w_lg_w_piso_sipo_q_range186w191w192w & wire_w_lg_w_lg_w_piso_sipo_q_range176w181w182w & wire_w_lg_w_lg_w_piso_sipo_q_range166w171w172w & wire_w_lg_w_lg_ufm_drdout160w161w);
	piso_sipo_q <= ( piso_sipo_dffe(15 DOWNTO 0));
	program1 <= program_dffe;
	q0 <= wire_cntr2_q(0);
	q1 <= wire_cntr2_q(1);
	q2 <= wire_cntr2_q(2);
	q3 <= wire_cntr2_q(3);
	q4 <= wire_cntr2_q(4);
	read_data_en <= (in_read_data_en AND read_op);
	read_drclk <= (in_read_drclk AND read_op);
	read_drshft <= (in_read_drshft AND read_op);
	read_op <= wire_w_lg_w_lg_w_lg_tmp_read36w37w38w(0);
	real_decode <= start_decode;
	shiftin <= ( A(7 DOWNTO 0) & "0");
	start_decode <= (wire_w_lg_ufm_bgpbusy25w(0) AND ((wire_w_lg_w_lg_w_lg_mux_nread20w21w22w(0) OR wire_w_lg_w_lg_mux_nread18w19w(0)) OR ((mux_nread AND mux_nwrite) AND wire_w_lg_mux_nerase14w(0))));
	start_op <= (hold_decode OR stop_op);
	stop_op <= ((((q4 AND q3) AND wire_w_lg_q253w(0)) AND q1) AND q0);
	tmp_add_en <= (wire_w_lg_q43w(0) AND wire_w_lg_w_lg_q363w64w(0));
	tmp_add_load <= (NOT (wire_w_lg_q43w(0) AND (((wire_w_lg_w_lg_q363w128w(0) OR wire_w_lg_w_lg_q363w127w(0)) OR wire_w_lg_w_lg_q363w126w(0)) OR (wire_w_lg_q3124w(0) AND wire_w_lg_q161w(0)))));
	tmp_arclk <= (gated1 AND wire_w_lg_ufm_osc321w(0));
	tmp_arclk0 <= (wire_w_lg_q43w(0) AND (wire_w_lg_q363w(0) OR (wire_w_lg_w_lg_q253w62w(0) AND wire_w_lg_q059w(0))));
	tmp_ardin <= A(8);
	tmp_arshft <= add_en;
	tmp_data_valid2 <= (stop_op AND read_op);
	tmp_decode <= ((wire_w_lg_w_lg_w_lg_tmp_read36w37w38w(0) OR wire_w_lg_w_lg_tmp_read34w35w(0)) OR ((tmp_read AND tmp_write) AND wire_w_lg_tmp_erase30w(0)));
	tmp_di <= ( datain(7 DOWNTO 0) & "00000001");
	tmp_drclk <= (gated2 AND wire_w_lg_ufm_osc321w(0));
	tmp_drdin <= piso_sipo_dffe(15);
	tmp_erase <= deco3_dffe;
	tmp_read <= deco1_dffe;
	tmp_write <= deco2_dffe;
	ufm_arclk <= tmp_arclk;
	ufm_ardin <= tmp_ardin;
	ufm_arshft <= tmp_arshft;
	ufm_bgpbusy <= wire_maxii_ufm_block1_bgpbusy;
	ufm_busy <= wire_maxii_ufm_block1_busy;
	ufm_drclk <= tmp_drclk;
	ufm_drdin <= tmp_drdin;
	ufm_drdout <= wire_maxii_ufm_block1_drdout;
	ufm_drshft <= drshft;
	ufm_erase <= ((erase OR ufm_busy) AND erase_op);
	ufm_osc <= wire_maxii_ufm_block1_osc;
	ufm_oscena <= oscena;
	ufm_program <= (in_program AND write_op);
	write_data_en <= (in_write_data_en AND write_op);
	write_data_load <= (in_write_data_load AND write_op);
	write_drclk <= (in_write_drclk AND write_op);
	write_drshft <= (in_write_drshft AND write_op);
	write_op <= wire_w_lg_w_lg_tmp_read34w35w(0);
	X_var <= wire_w_lg_shiftin143w;
	Y_var <= wire_w_lg_addr144w;
	Z_var <= (X_var OR Y_var);
	wire_w_piso_sipo_q_range166w(0) <= piso_sipo_q(0);
	wire_w_piso_sipo_q_range266w(0) <= piso_sipo_q(10);
	wire_w_piso_sipo_q_range276w(0) <= piso_sipo_q(11);
	wire_w_piso_sipo_q_range286w(0) <= piso_sipo_q(12);
	wire_w_piso_sipo_q_range296w(0) <= piso_sipo_q(13);
	wire_w_piso_sipo_q_range306w(0) <= piso_sipo_q(14);
	wire_w_piso_sipo_q_range176w(0) <= piso_sipo_q(1);
	wire_w_piso_sipo_q_range186w(0) <= piso_sipo_q(2);
	wire_w_piso_sipo_q_range196w(0) <= piso_sipo_q(3);
	wire_w_piso_sipo_q_range206w(0) <= piso_sipo_q(4);
	wire_w_piso_sipo_q_range216w(0) <= piso_sipo_q(5);
	wire_w_piso_sipo_q_range226w(0) <= piso_sipo_q(6);
	wire_w_piso_sipo_q_range236w(0) <= piso_sipo_q(7);
	wire_w_piso_sipo_q_range246w(0) <= piso_sipo_q(8);
	wire_w_piso_sipo_q_range256w(0) <= piso_sipo_q(9);
	wire_w_tmp_di_range156w(0) <= tmp_di(0);
	wire_w_tmp_di_range258w(0) <= tmp_di(10);
	wire_w_tmp_di_range268w(0) <= tmp_di(11);
	wire_w_tmp_di_range278w(0) <= tmp_di(12);
	wire_w_tmp_di_range288w(0) <= tmp_di(13);
	wire_w_tmp_di_range298w(0) <= tmp_di(14);
	wire_w_tmp_di_range308w(0) <= tmp_di(15);
	wire_w_tmp_di_range168w(0) <= tmp_di(1);
	wire_w_tmp_di_range178w(0) <= tmp_di(2);
	wire_w_tmp_di_range188w(0) <= tmp_di(3);
	wire_w_tmp_di_range198w(0) <= tmp_di(4);
	wire_w_tmp_di_range208w(0) <= tmp_di(5);
	wire_w_tmp_di_range218w(0) <= tmp_di(6);
	wire_w_tmp_di_range228w(0) <= tmp_di(7);
	wire_w_tmp_di_range238w(0) <= tmp_di(8);
	wire_w_tmp_di_range248w(0) <= tmp_di(9);
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (add_en = '1') THEN A <= ( Z_var);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN data_valid_out_reg <= wire_data_valid_reg_w_lg_q100w(0);
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (data_valid_en = '1') THEN data_valid_reg <= tmp_data_valid2;
			END IF;
		END IF;
	END PROCESS;
	wire_data_valid_reg_w_lg_q100w(0) <= data_valid_reg AND wire_w_lg_tmp_decode99w(0);
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (start_op = '1') THEN deco1_dffe <= mux_nread;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (start_op = '1') THEN deco2_dffe <= mux_nwrite;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (start_op = '1') THEN deco3_dffe <= mux_nerase;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN decode_dffe <= copy_tmp_decode;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN gated_clk1_dffe <= busy_arclk;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN gated_clk2_dffe <= busy_drclk;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (data_en = '1') THEN piso_sipo_dffe <= ( piso_sipo_d(15 DOWNTO 0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_busy, wire_program_dffe_clrn)
	BEGIN
		IF (wire_program_dffe_clrn = '0') THEN program_dffe <= '0';
		ELSIF (ufm_busy = '0' AND ufm_busy'event) THEN program_dffe <= (ufm_program OR ufm_erase);
		END IF;
	END PROCESS;
	wire_program_dffe_clrn <= (NOT (stop_op OR ((((wire_w_lg_q43w(0) AND wire_w_lg_q363w(0)) AND wire_w_lg_q253w(0)) AND wire_w_lg_q161w(0)) AND wire_w_lg_q059w(0))));
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN real_decode2_dffe <= real_decode_dffe;
		END IF;
	END PROCESS;
	wire_real_decode2_dffe_w_lg_q27w(0) <= NOT real_decode2_dffe;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN real_decode_dffe <= start_decode;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(0) = '1') THEN tmp_do(0) <= wire_tmp_do_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(1) = '1') THEN tmp_do(1) <= wire_tmp_do_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(2) = '1') THEN tmp_do(2) <= wire_tmp_do_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(3) = '1') THEN tmp_do(3) <= wire_tmp_do_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(4) = '1') THEN tmp_do(4) <= wire_tmp_do_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(5) = '1') THEN tmp_do(5) <= wire_tmp_do_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(6) = '1') THEN tmp_do(6) <= wire_tmp_do_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(7) = '1') THEN tmp_do(7) <= wire_tmp_do_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_tmp_do_d <= ( piso_sipo_q(15 DOWNTO 8));
	loop2 : FOR i IN 0 TO 7 GENERATE
		wire_tmp_do_ena(i) <= wire_data_valid_reg_w_lg_q100w(0);
	END GENERATE loop2;
	wire_cntr2_cnt_en <= wire_w_lg_w_lg_w_lg_ufm_program45w46w47w(0);
	wire_w_lg_w_lg_w_lg_ufm_program45w46w47w(0) <= (NOT (ufm_program OR ufm_erase)) OR program1;
	cntr2 :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_modulus => 28,
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 5
	  )
	  PORT MAP ( 
		clk_en => tmp_decode,
		clock => ufm_osc,
		cnt_en => wire_cntr2_cnt_en,
		q => wire_cntr2_q
	  );
	maxii_ufm_block1 :  maxii_ufm
	  GENERIC MAP (
		ADDRESS_WIDTH => 9,
		ERASE_TIME => 500000000,
		INIT_FILE => "tstdata.mif",
		mem1 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001000011111111000011111111111100001110111111110000110111111111000011001111111100001011111111110000101011111111000010011111111100001000111111110000011111111111000001101111111100000101111111110000010011111111000000111111111100000010111111110000000111111111",
		mem10 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem11 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem12 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem13 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem14 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem15 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem16 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem2 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem3 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem4 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem5 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem6 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem7 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem8 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem9 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		OSC_SIM_SETTING => 180000,
		PROGRAM_TIME => 1600000
	  )
	  PORT MAP ( 
		arclk => ufm_arclk,
		ardin => ufm_ardin,
		arshft => ufm_arshft,
		bgpbusy => wire_maxii_ufm_block1_bgpbusy,
		busy => wire_maxii_ufm_block1_busy,
		drclk => ufm_drclk,
		drdin => ufm_drdin,
		drdout => wire_maxii_ufm_block1_drdout,
		drshft => ufm_drshft,
		erase => ufm_erase,
		osc => wire_maxii_ufm_block1_osc,
		oscena => ufm_oscena,
		program => ufm_program
	  );

 END RTL; --flash_altufm_parallel_22p
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY flash IS
	PORT
	(
		addr		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		datain		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		nerase		: IN STD_LOGIC ;
		nread		: IN STD_LOGIC ;
		nwrite		: IN STD_LOGIC ;
		data_valid		: OUT STD_LOGIC ;
		dataout		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		nbusy		: OUT STD_LOGIC 
	);
END flash;


ARCHITECTURE RTL OF flash IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "altufm_parallel";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "access_mode=READ_WRITE;erase_time=500000000;intended_device_family=MAX II;lpm_file=tstdata.mif;osc_frequency=180000;program_time=1600000;width_address=9;width_data=8;width_ufm_address=9;";
	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC ;
	SIGNAL sub_wire2	: STD_LOGIC ;



	COMPONENT flash_altufm_parallel_22p
	PORT (
			dataout	: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			addr	: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
			datain	: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			nwrite	: IN STD_LOGIC ;
			nerase	: IN STD_LOGIC ;
			data_valid	: OUT STD_LOGIC ;
			nread	: IN STD_LOGIC ;
			nbusy	: OUT STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	dataout    <= sub_wire0(7 DOWNTO 0);
	data_valid    <= sub_wire1;
	nbusy    <= sub_wire2;

	flash_altufm_parallel_22p_component : flash_altufm_parallel_22p
	PORT MAP (
		addr => addr,
		datain => datain,
		nwrite => nwrite,
		nerase => nerase,
		nread => nread,
		dataout => sub_wire0,
		data_valid => sub_wire1,
		nbusy => sub_wire2
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "MAX II"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_PART STRING ""
-- Retrieval info: PRIVATE: INTERFACE_CHOICE NUMERIC "1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: VERSION_NUMBER NUMERIC "0"
-- Retrieval info: CONSTANT: ACCESS_MODE STRING "READ_WRITE"
-- Retrieval info: CONSTANT: ERASE_TIME NUMERIC "500000000"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "MAX II"
-- Retrieval info: CONSTANT: LPM_FILE STRING "tstdata.mif"
-- Retrieval info: CONSTANT: OSC_FREQUENCY NUMERIC "180000"
-- Retrieval info: CONSTANT: PROGRAM_TIME NUMERIC "1600000"
-- Retrieval info: CONSTANT: WIDTH_ADDRESS NUMERIC "9"
-- Retrieval info: CONSTANT: WIDTH_DATA NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_UFM_ADDRESS NUMERIC "9"
-- Retrieval info: USED_PORT: addr 0 0 9 0 INPUT NODEFVAL addr[8..0]
-- Retrieval info: USED_PORT: data_valid 0 0 0 0 OUTPUT NODEFVAL data_valid
-- Retrieval info: USED_PORT: datain 0 0 8 0 INPUT NODEFVAL datain[7..0]
-- Retrieval info: USED_PORT: dataout 0 0 8 0 OUTPUT NODEFVAL dataout[7..0]
-- Retrieval info: USED_PORT: nbusy 0 0 0 0 OUTPUT NODEFVAL nbusy
-- Retrieval info: USED_PORT: nerase 0 0 0 0 INPUT NODEFVAL nerase
-- Retrieval info: USED_PORT: nread 0 0 0 0 INPUT NODEFVAL nread
-- Retrieval info: USED_PORT: nwrite 0 0 0 0 INPUT NODEFVAL nwrite
-- Retrieval info: CONNECT: @nwrite 0 0 0 0 nwrite 0 0 0 0
-- Retrieval info: CONNECT: @nerase 0 0 0 0 nerase 0 0 0 0
-- Retrieval info: CONNECT: @datain 0 0 8 0 datain 0 0 8 0
-- Retrieval info: CONNECT: @nread 0 0 0 0 nread 0 0 0 0
-- Retrieval info: CONNECT: @addr 0 0 9 0 addr 0 0 9 0
-- Retrieval info: CONNECT: nbusy 0 0 0 0 @nbusy 0 0 0 0
-- Retrieval info: CONNECT: data_valid 0 0 0 0 @data_valid 0 0 0 0
-- Retrieval info: CONNECT: dataout 0 0 8 0 @dataout 0 0 8 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL flash.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL flash.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL flash.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL flash.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL flash_inst.vhd TRUE
-- Retrieval info: LIB_FILE: lpm
-- Retrieval info: LIB_FILE: maxii
